module segment7(input logic clk, input logic [3:0] s, output logic [2:0] led, output logic [6:0] seg);

always_comb begin :
    case (s)
        4'hf: seg = 7'b0001110;
        4'he: seg = 7'b0000110;
        4'hd: seg = 7'b0110000;
        4'hc: seg = 7'b1001100;
        4'hb: seg = 7'b0011000;
        4'ha: seg = 7'b0000010;
        4'h9: seg = 7'b0000001;
        4'h8: seg = 7'b0000000;
        4'h7: seg = 7'b1100011;
        4'h6: seg = 7'b0001000;
        4'h5: seg = 7'b0001001;
        4'h4: seg = 7'b0010011;
        4'h3: seg = 7'b0100001;
        4'h2: seg = 7'b0100100;
        4'h1: seg = 7'b1110011;
        4'h0: seg = 7'b1000000;   
        default: seg = 7'b1111111;
    endcase
    end
endmodule
